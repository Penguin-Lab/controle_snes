library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity mario_sprite is
    Port ( clock : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           trigger : in  STD_LOGIC;
           hc : in  INTEGER;
           vc : in  INTEGER;
			  Ax : in  STD_LOGIC_VECTOR (7 downto 0);
			  B  : in  STD_LOGIC;
           mario_on : out  STD_LOGIC;
           rm : out  STD_LOGIC_VECTOR (2 downto 0);
           gm : out  STD_LOGIC_VECTOR (2 downto 0);
           bm : out  STD_LOGIC_VECTOR (1 downto 0));
end mario_sprite;

architecture Behavioral of mario_sprite is

signal hm : integer := 192;
signal vm : integer := 468;
signal Ax_digital : integer;
signal marrom, vermelho, rosa : std_logic;
signal direction : std_logic := '0';
type mario_bits is array (0 to 31) of std_logic_vector (0 to 31);
signal vermelho_bits,rosa_bits,marrom_bits : mario_bits;
signal index_h, index_v : integer range 0 to 31;
signal sprite : integer := 0;
signal pulo : std_logic := '0';
signal estado_pulo,prox_estado : integer := 0;
constant altura : integer := 64;

begin

-- FSM pulo
process(clock,reset)
begin
if reset = '1' then
	vm <= 468;
	estado_pulo <= 0;
elsif rising_edge(clock) then
	if trigger = '1' then
		estado_pulo <= prox_estado;
		if estado_pulo = 1 then
			vm <= vm - 16;
			if vm <= (468-altura) then
				vm <= (468-altura);
			end if;
		elsif estado_pulo = 2 then
			vm <= vm + 16;
			if vm >= 468 then
				vm <= 468;
			end if;
		end if;
	end if;
end if;
end process;

process(B,vm,estado_pulo)
begin
	case estado_pulo is
	when 0 =>
		if B = '1' then
			prox_estado <= 1;
		else
			prox_estado <= 0;
		end if;
	when 1 =>
		if vm <= (468-altura) then
			prox_estado <= 2;
		else
			prox_estado <= 1;
		end if;
	when others =>
		if vm = 468 then
			prox_estado <= 0;
		else
			prox_estado <= 2;
		end if;
	end case;
end process;

pulo <= '0' when estado_pulo = 0 else
		  '1';

-- FSM sprites

process(clock,reset)
begin
if reset = '1' then
	sprite <= 0;
elsif rising_edge(clock) then
	if trigger = '1' then
		if pulo = '1' then
			sprite <= 4;
		elsif pulo = '0' and ((Ax_digital > 140 and hm < (799-32)) or (Ax_digital < 115 and hm > (160+32))) then
			sprite <= sprite + 1;
			if sprite >= 3 then
				sprite <= 1;
			end if;
		else
			sprite <= 0;
		end if;
	end if;
end if;
end process;

Ax_digital <= 255 - to_integer(unsigned(Ax));

process(clock, reset)
begin
if reset = '1' then
	hm <= 192;
	direction <= '0';
elsif rising_edge(clock) then
	if trigger = '1' then
		if Ax_digital > 140 and hm < (799-32) then
			hm <= hm + 10;
			direction <= '0';
		elsif Ax_digital < 115 and hm > (160+32) then
			hm <= hm - 10;
			direction <= '1';
		end if;
	end if;
end if;
end process;

-- Cores
index_h <= (hc - hm) when direction = '0' and (hc >= hm and hc < (hm+32)) else
			(31 - hc + hm) when direction = '1' and (hc >= hm and hc < (hm+32)) else
			0;
index_v <= (vc - vm) when (vc >= vm and vc < (vm+32)) else
			0;

process(hc,hm,vc,vm)
begin
if (hc >= hm and hc < (hm+32)) and (vc >= vm and vc < (vm+32)) then
	vermelho <= vermelho_bits(index_v)(index_h);
	rosa <= rosa_bits(index_v)(index_h);
	marrom <= marrom_bits(index_v)(index_h);
else
	vermelho <= '0';
	rosa <= '0';
	marrom <= '0';
end if;
end process;

-- Saidas
mario_on <= '1' when vermelho = '1' or rosa = '1' or marrom = '1' else '0';

rm <= "101" when vermelho = '1' else
		"111" when rosa = '1' else
		"010" when marrom = '1' else
		"000";
gm <= "000" when vermelho = '1' else
		"110" when rosa = '1' else
		"001" when marrom = '1' else
		"000";
bm <= "00" when vermelho = '1' else
		"10" when rosa = '1' else
		"00" when marrom = '1' else
		"00";

-- Mario bits
-- Sprite parado (0)
-- Sprite andando1 (1)
-- Sprite andando2 (2)
-- Sprite andando3 (3)
-- Sprite pulando (4)
vermelho_bits <= (
			"00000000001111111111000000000000",
			"00000000001111111111000000000000",
			"00000000111111111111111111000000",
			"00000000111111111111111111000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000011000000000000000000",
			"00000000000011000000000000000000",
			"00000000000011000011000000000000",
			"00000000000011000011000000000000",
			"00000000000011111111000000000000",
			"00000000000011111111000000000000",
			"00000000001100111100110000000000",
			"00000000001100111100110000000000",
			"00000000001111111111110000000000",
			"00000000001111111111110000000000",
			"00000000111111111111111100000000",
			"00000000111111111111111100000000",
			"00000000111111000011111100000000",
			"00000000111111000011111100000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			) when sprite = 0 else
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000011111111110000000000",
			"00000000000011111111110000000000",
			"00000000001111111111111111110000",
			"00000000001111111111111111110000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000011000000000000",
			"00000000000000000011000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000001100000000000000000000",
			"00000000001100000000000000000000",
			"00000000001111111111111100000000",
			"00000000001111111111111100000000",
			"00000000111111111111111100000000",
			"00000000111111111111111100000000",
			"00000000111111001111110000000000",
			"00000000111111001111110000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			) when sprite = 1 else
			(
			"00000000001111111111000000000000",
			"00000000001111111111000000000000",
			"00000000111111111111111111000000",
			"00000000111111111111111111000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000011000000000000000000",
			"00000000000011000000000000000000",
			"00000000000000111100000000000000",
			"00000000000000111100000000000000",
			"00000000000011110011110000000000",
			"00000000000011110011110000000000",
			"00000000000000111111111100000000",
			"00000000000000111111111100000000",
			"00000011000000000011111100000000",
			"00000011000000000011111100000000",
			"00000000110000001111110000000000",
			"00000000110000001111110000000000",
			"00000000001111110000000000000000",
			"00000000001111110000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			) when sprite = 2 else
			(
			"00000000001111111111000000000000",
			"00000000001111111111000000000000",
			"00000000111111111111111111000000",
			"00000000111111111111111111000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000011110000000000000000",
			"00000000000011110000000000000000",
			"00000000000011111100000000000000",
			"00000000000011111100000000000000",
			"00000000000011001111110000000000",
			"00000000000011001111110000000000",
			"00000000111111111111110000000000",
			"00000000111111111111110000000000",
			"00000011111111111111111100000000",
			"00000011111111111111111100000000",
			"00001111111111111111111100000000",
			"00001111111111111111111100000000",
			"00000011111100000011111100000000",
			"00000011111100000011111100000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			) when sprite = 3 else
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000011111111110000000000",
			"00000000000011111111110000000000",
			"00000000001111111111111111110000",
			"00000000001111111111111111110000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000110000001100000000",
			"00000000000000110000001100000000",
			"00000000000000001100000011000000",
			"00000000000000001100000011000000",
			"00000000000000001111111111000000",
			"00000000000000001111111111000000",
			"00000000111100111100111100110000",
			"00000000111100111100111100110000",
			"00000000111111111111111111110000",
			"00000000111111111111111111110000",
			"00000000001111111111111111110000",
			"00000000001111111111111111110000",
			"00000000111111111111110000000000",
			"00000000111111111111110000000000",
			"00000000111111110000000000000000",
			"00000000111111110000000000000000"
			);

rosa_bits <= (
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000111100110000000000",
			"00000000000000111100110000000000",
			"00000000110011111100111111000000",
			"00000000110011111100111111000000",
			"00000000110000111111001111110000",
			"00000000110000111111001111110000",
			"00000000001111111100000000000000",
			"00000000001111111100000000000000",
			"00000000001111111111111100000000",
			"00000000001111111111111100000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00001111000011000011000011110000",
			"00001111000011000011000011110000",
			"00001111110000000000001111110000",
			"00001111110000000000001111110000",
			"00001111000000000000000011110000",
			"00001111000000000000000011110000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			) when sprite = 0 else
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000001111001100000000",
			"00000000000000001111001100000000",
			"00000000001100111111001111110000",
			"00000000001100111111001111110000",
			"00000000001100001111110011110000",
			"00000000001100001111110011110000",
			"00000000000011111111000000000000",
			"00000000000011111111000000000000",
			"00000000000011111111111111000000",
			"00000000000011111111111111000000",
			"00000000000000000000000011000000",
			"00000000000000000000000011000000",
			"00000000110000000000001111110000",
			"00000000110000000000001111110000",
			"00000011110000000000001111000000",
			"00000011110000000000001111000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			) when sprite = 1 else
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000111100110000000000",
			"00000000000000111100110000000000",
			"00000000110011111100111111000000",
			"00000000110011111100111111000000",
			"00000000110000111111001111110000",
			"00000000110000111111001111110000",
			"00000000001111111100000000000000",
			"00000000001111111100000000000000",
			"00000000001111111111111100000000",
			"00000000001111111111111100000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000001100001100000000",
			"00000000000000001100001100000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000011111100000000000000",
			"00000000000011111100000000000000",
			"00000000000011110000000000000000",
			"00000000000011110000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			) when sprite = 2 else
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000111100110000000000",
			"00000000000000111100110000000000",
			"00000000110011111100111111000000",
			"00000000110011111100111111000000",
			"00000000110000111111001111110000",
			"00000000110000111111001111110000",
			"00000000001111111100000000000000",
			"00000000001111111100000000000000",
			"00000000001111111111111100000000",
			"00000000001111111111111100000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"11110000000000000000000011111100",
			"11110000000000000000000011111100",
			"11111100000000110000000000111100",
			"11111100000000110000000000111100",
			"11110000000000000000000000000000",
			"11110000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			) when sprite = 3 else
			(
			"00000000000000000000000000111111",
			"00000000000000000000000000111111",
			"00000000000000000000000000111111",
			"00000000000000000000000000111111",
			"00000000000000000000000000001111",
			"00000000000000000000000000001111",
			"00000000000000001111001100000000",
			"00000000000000001111001100000000",
			"00000000001100111111001111000000",
			"00000000001100111111001111000000",
			"00000000001100001111110011111100",
			"00000000001100001111110011111100",
			"00000000000011111111000000000000",
			"00000000000011111111000000000000",
			"00000000000011111111111111000000",
			"00000000000011111111111111000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"11110000000000000000000000000000",
			"11110000000000000000000000000000",
			"11111100000000000011000011000000",
			"11111100000000000011000011000000",
			"00110000000000000000000000000000",
			"00110000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000"
			);

marrom_bits <= 
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000111111000011000000000000",
			"00000000111111000011000000000000",
			"00000011001100000011000000000000",
			"00000011001100000011000000000000",
			"00000011001111000000110000000000",
			"00000011001111000000110000000000",
			"00000011110000000011111111000000",
			"00000011110000000011111111000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000111100111111000000000000",
			"00000000111100111111000000000000",
			"00000011111100111100111111000000",
			"00000011111100111100111111000000",
			"00001111111100000000111111110000",
			"00001111111100000000111111110000",
			"00000000110000000000001100000000",
			"00000000110000000000001100000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000011111100000000111111000000",
			"00000011111100000000111111000000",
			"00001111111100000000111111110000",
			"00001111111100000000111111110000"
			) when sprite = 0 else
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000001111110000110000000000",
			"00000000001111110000110000000000",
			"00000000110011000000110000000000",
			"00000000110011000000110000000000",
			"00000000110011110000001100000000",
			"00000000110011110000001100000000",
			"00000000111100000000111111110000",
			"00000000111100000000111111110000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000001111111100110000000000",
			"00000000001111111100110000000000",
			"00000000001111111111110000000000",
			"00000000001111111111110000000000",
			"00000000000011111111110000000000",
			"00000000000011111111110000000000",
			"00000011110000000000000000000000",
			"00000011110000000000000000000000",
			"00000011000000000000000000000000",
			"00000011000000000000000000000000",
			"00001111000000000000000000000000",
			"00001111000000000000000000000000",
			"00001100000000111111000000000000",
			"00001100000000111111000000000000",
			"00000000000000111111110000000000",
			"00000000000000111111110000000000"
			) when sprite = 1 else
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000111111000011000000000000",
			"00000000111111000011000000000000",
			"00000011001100000011000000000000",
			"00000011001100000011000000000000",
			"00000011001111000000110000000000",
			"00000011001111000000110000000000",
			"00000011110000000011111111000000",
			"00000011110000000011111111000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000111100111111000000000000",
			"00000000111100111111000000000000",
			"00000011111111000011110000000000",
			"00000011111111000011110000000000",
			"00000011111100000000000000000000",
			"00000011111100000000000000000000",
			"00000011111111000000000000000000",
			"00000011111111000000000000000000",
			"00000000111100000000000000000000",
			"00000000111100000000000000000000",
			"00000000001100000000000000000000",
			"00000000001100000000000000000000",
			"00000000000000001111110000000000",
			"00000000000000001111110000000000",
			"00000000001111111111111100000000",
			"00000000001111111111111100000000",
			"00000000001111111100000000000000",
			"00000000001111111100000000000000"
			) when sprite = 2 else
			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000111111000011000000000000",
			"00000000111111000011000000000000",
			"00000011001100000011000000000000",
			"00000011001100000011000000000000",
			"00000011001111000000110000000000",
			"00000011001111000000110000000000",
			"00000011110000000011111111000000",
			"00000011110000000011111111000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00001111111100001111000000000000",
			"00001111111100001111000000000000",
			"00001111111100000011111100000000",
			"00001111111100000011111100000000",
			"00000000111100000000001111000000",
			"00000000111100000000001111000000",
			"00000000000000000000000000110000",
			"00000000000000000000000000110000",
			"00000000000000000000000011110000",
			"00000000000000000000000011110000",
			"00000000000000000000000011110000",
			"00000000000000000000000011110000",
			"00111100000000000000000011110000",
			"00111100000000000000000011110000",
			"00111111000000000000000000000000",
			"00111111000000000000000000000000",
			"00001111110000000000000000000000",
			"00001111110000000000000000000000"
			) when sprite = 3 else

			(
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000000000000000000000000000",
			"00000000001111110000110000111111",
			"00000000001111110000110000111111",
			"00000000110011000000110000111111",
			"00000000110011000000110000111111",
			"00000000110011110000001100000011",
			"00000000110011110000001100000011",
			"00000000111100000000111111111100",
			"00000000111100000000111111111100",
			"00000000000000000000000000110000",
			"00000000000000000000000000110000",
			"00001111111111001111110011000000",
			"00001111111111001111110011000000",
			"00111111111111110011111100000011",
			"00111111111111110011111100000011",
			"00001111111111110000000000000011",
			"00001111111111110000000000000011",
			"00000000000011000000000000001111",
			"00000000000011000000000000001111",
			"00000011000000000000000000001111",
			"00000011000000000000000000001111",
			"00001111110000000000000000001111",
			"00001111110000000000000000001111",
			"00111111000000000000000000000000",
			"00111111000000000000000000000000",
			"00110000000000000000000000000000",
			"00110000000000000000000000000000"
			);

end Behavioral;

